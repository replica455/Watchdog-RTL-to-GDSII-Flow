magic
tech scmos
timestamp 1656334919
<< metal1 >>
rect 280 303 282 307
rect 286 303 289 307
rect 293 303 296 307
rect 210 278 217 281
rect 142 268 153 271
rect 166 268 190 271
rect 234 268 257 271
rect 270 268 297 271
rect 114 258 121 261
rect 104 203 106 207
rect 110 203 113 207
rect 117 203 120 207
rect 286 188 294 191
rect 38 148 54 151
rect 150 148 158 151
rect 138 138 145 141
rect 126 128 137 131
rect 94 118 102 121
rect 250 118 251 122
rect 280 103 282 107
rect 286 103 289 107
rect 293 103 296 107
rect 14 78 25 81
rect 110 78 118 81
rect 14 68 22 71
rect 78 68 89 71
rect 106 68 142 71
rect 182 68 190 71
rect 222 68 230 71
rect 246 68 270 71
rect 286 68 313 71
rect 122 58 134 61
rect 346 58 353 61
rect 358 58 377 61
rect 406 38 414 41
rect 104 3 106 7
rect 110 3 113 7
rect 117 3 120 7
<< m2contact >>
rect 282 303 286 307
rect 289 303 293 307
rect 174 278 178 282
rect 198 278 202 282
rect 206 278 210 282
rect 246 278 250 282
rect 134 266 138 270
rect 190 268 194 272
rect 230 268 234 272
rect 350 268 354 272
rect 38 258 42 262
rect 62 258 66 262
rect 110 258 114 262
rect 182 258 186 262
rect 222 258 226 262
rect 238 258 242 262
rect 302 258 306 262
rect 318 258 322 262
rect 358 258 362 262
rect 94 218 98 222
rect 414 218 418 222
rect 106 203 110 207
rect 113 203 117 207
rect 166 188 170 192
rect 294 188 298 192
rect 222 168 226 172
rect 206 158 210 162
rect 254 158 258 162
rect 54 148 58 152
rect 62 148 66 152
rect 158 148 162 152
rect 190 148 194 152
rect 214 148 218 152
rect 270 148 274 152
rect 334 147 338 151
rect 134 138 138 142
rect 198 138 202 142
rect 238 138 242 142
rect 262 138 266 142
rect 350 138 354 142
rect 118 128 122 132
rect 158 128 162 132
rect 222 128 226 132
rect 102 118 106 122
rect 174 118 178 122
rect 246 118 250 122
rect 398 118 402 122
rect 282 103 286 107
rect 289 103 293 107
rect 54 88 58 92
rect 174 88 178 92
rect 334 88 338 92
rect 6 78 10 82
rect 118 78 122 82
rect 150 78 154 82
rect 158 78 162 82
rect 166 78 170 82
rect 230 78 234 82
rect 262 78 266 82
rect 342 78 346 82
rect 22 68 26 72
rect 30 68 34 72
rect 102 68 106 72
rect 142 68 146 72
rect 190 68 194 72
rect 214 66 218 70
rect 230 68 234 72
rect 270 68 274 72
rect 382 68 386 72
rect 46 58 50 62
rect 70 58 74 62
rect 118 58 122 62
rect 134 58 138 62
rect 190 58 194 62
rect 198 58 202 62
rect 238 58 242 62
rect 254 58 258 62
rect 318 58 322 62
rect 342 58 346 62
rect 390 58 394 62
rect 366 48 370 52
rect 414 38 418 42
rect 106 3 110 7
rect 113 3 117 7
<< metal2 >>
rect 280 303 282 307
rect 286 303 289 307
rect 293 303 296 307
rect 198 282 201 288
rect 166 278 174 281
rect 238 278 246 281
rect 134 270 137 278
rect 42 258 46 261
rect 106 258 110 261
rect 62 162 65 258
rect 62 152 65 158
rect 54 92 57 148
rect 94 142 97 218
rect 104 203 106 207
rect 110 203 113 207
rect 117 203 120 207
rect 166 192 169 278
rect 174 261 177 278
rect 194 268 201 271
rect 174 258 182 261
rect 190 152 193 168
rect 118 132 121 138
rect 6 72 9 78
rect 18 68 22 71
rect 30 52 33 68
rect 70 62 73 78
rect 102 72 105 118
rect 118 62 121 78
rect 134 62 137 138
rect 158 132 161 148
rect 198 142 201 268
rect 206 222 209 278
rect 218 258 222 261
rect 230 172 233 268
rect 238 262 241 278
rect 298 258 302 261
rect 238 192 241 258
rect 318 252 321 258
rect 290 188 294 191
rect 226 168 230 171
rect 194 138 198 141
rect 162 128 166 131
rect 174 112 177 118
rect 142 72 145 98
rect 206 92 209 158
rect 214 122 217 148
rect 254 142 257 158
rect 350 152 353 268
rect 358 252 361 258
rect 382 152 385 168
rect 414 152 417 218
rect 226 128 230 131
rect 178 88 182 91
rect 150 82 153 88
rect 158 62 161 78
rect 166 72 169 78
rect 194 68 201 71
rect 198 62 201 68
rect 214 70 217 118
rect 238 102 241 138
rect 226 78 230 81
rect 238 71 241 98
rect 246 82 249 118
rect 262 92 265 138
rect 270 122 273 148
rect 234 68 241 71
rect 254 62 257 88
rect 262 82 265 88
rect 270 72 273 118
rect 280 103 282 107
rect 286 103 289 107
rect 293 103 296 107
rect 334 92 337 147
rect 350 142 353 148
rect 338 78 342 81
rect 50 58 54 61
rect 186 58 190 61
rect 234 58 238 61
rect 314 58 318 61
rect 346 58 350 61
rect 366 52 369 118
rect 382 72 385 148
rect 394 118 398 121
rect 386 58 390 61
rect 414 42 417 48
rect 104 3 106 7
rect 110 3 113 7
rect 117 3 120 7
<< m3contact >>
rect 282 303 286 307
rect 289 303 293 307
rect 198 288 202 292
rect 134 278 138 282
rect 46 258 50 262
rect 102 258 106 262
rect 62 158 66 162
rect 106 203 110 207
rect 113 203 117 207
rect 190 168 194 172
rect 94 138 98 142
rect 118 138 122 142
rect 70 78 74 82
rect 6 68 10 72
rect 14 68 18 72
rect 214 258 218 262
rect 206 218 210 222
rect 294 258 298 262
rect 318 248 322 252
rect 238 188 242 192
rect 286 188 290 192
rect 230 168 234 172
rect 190 138 194 142
rect 166 128 170 132
rect 174 108 178 112
rect 142 98 146 102
rect 358 248 362 252
rect 382 168 386 172
rect 254 138 258 142
rect 230 128 234 132
rect 214 118 218 122
rect 150 88 154 92
rect 182 88 186 92
rect 206 88 210 92
rect 158 78 162 82
rect 166 68 170 72
rect 238 98 242 102
rect 222 78 226 82
rect 350 148 354 152
rect 382 148 386 152
rect 414 148 418 152
rect 270 118 274 122
rect 254 88 258 92
rect 262 88 266 92
rect 246 78 250 82
rect 282 103 286 107
rect 289 103 293 107
rect 366 118 370 122
rect 334 78 338 82
rect 54 58 58 62
rect 158 58 162 62
rect 182 58 186 62
rect 230 58 234 62
rect 310 58 314 62
rect 350 58 354 62
rect 390 118 394 122
rect 382 58 386 62
rect 30 48 34 52
rect 414 48 418 52
rect 106 3 110 7
rect 113 3 117 7
<< metal3 >>
rect 280 303 282 307
rect 286 303 289 307
rect 294 303 296 307
rect 198 281 201 288
rect 138 278 201 281
rect 50 258 102 261
rect 218 258 294 261
rect 318 258 361 261
rect 318 252 321 258
rect 358 252 361 258
rect 206 212 209 218
rect 104 203 106 207
rect 110 203 113 207
rect 118 203 120 207
rect 242 188 286 191
rect 194 168 230 171
rect 234 168 382 171
rect -26 151 -22 152
rect 62 151 65 158
rect -26 148 350 151
rect 386 148 414 151
rect 98 138 118 141
rect 122 138 190 141
rect 194 138 254 141
rect 170 128 230 131
rect 218 118 270 121
rect 274 118 366 121
rect 370 118 390 121
rect 178 108 190 111
rect 280 103 282 107
rect 286 103 289 107
rect 294 103 296 107
rect 146 98 238 101
rect 174 88 182 91
rect 186 88 206 91
rect 210 88 254 91
rect 258 88 262 91
rect 150 81 153 88
rect 74 78 153 81
rect 162 78 206 81
rect 210 78 222 81
rect 250 78 334 81
rect -26 71 -22 72
rect -26 68 6 71
rect 18 68 166 71
rect 46 58 54 61
rect 58 58 158 61
rect 186 58 190 61
rect 234 58 310 61
rect 354 58 382 61
rect -26 51 -22 52
rect -26 48 30 51
rect 446 51 450 52
rect 418 48 450 51
rect 104 3 106 7
rect 110 3 113 7
rect 118 3 120 7
<< m4contact >>
rect 282 303 286 307
rect 290 303 293 307
rect 293 303 294 307
rect 206 208 210 212
rect 106 203 110 207
rect 114 203 117 207
rect 117 203 118 207
rect 190 108 194 112
rect 282 103 286 107
rect 290 103 293 107
rect 293 103 294 107
rect 206 78 210 82
rect 190 58 194 62
rect 106 3 110 7
rect 114 3 117 7
rect 117 3 118 7
<< metal4 >>
rect 280 303 282 307
rect 286 303 289 307
rect 294 303 296 307
rect 104 203 106 207
rect 110 203 113 207
rect 118 203 120 207
rect 190 62 193 108
rect 206 82 209 208
rect 280 103 282 107
rect 286 103 289 107
rect 294 103 296 107
rect 104 3 106 7
rect 110 3 113 7
rect 118 3 120 7
<< m5contact >>
rect 282 303 286 307
rect 289 303 290 307
rect 290 303 293 307
rect 106 203 110 207
rect 113 203 114 207
rect 114 203 117 207
rect 282 103 286 107
rect 289 103 290 107
rect 290 103 293 107
rect 106 3 110 7
rect 113 3 114 7
rect 114 3 117 7
<< metal5 >>
rect 286 303 289 307
rect 285 302 290 303
rect 295 302 296 307
rect 110 203 113 207
rect 109 202 114 203
rect 119 202 120 207
rect 286 103 289 107
rect 285 102 290 103
rect 295 102 296 107
rect 110 3 113 7
rect 109 2 114 3
rect 119 2 120 7
<< m6contact >>
rect 280 303 282 307
rect 282 303 285 307
rect 290 303 293 307
rect 293 303 295 307
rect 280 302 285 303
rect 290 302 295 303
rect 104 203 106 207
rect 106 203 109 207
rect 114 203 117 207
rect 117 203 119 207
rect 104 202 109 203
rect 114 202 119 203
rect 280 103 282 107
rect 282 103 285 107
rect 290 103 293 107
rect 293 103 295 107
rect 280 102 285 103
rect 290 102 295 103
rect 104 3 106 7
rect 106 3 109 7
rect 114 3 117 7
rect 117 3 119 7
rect 104 2 109 3
rect 114 2 119 3
<< metal6 >>
rect 104 207 120 310
rect 109 202 114 207
rect 119 202 120 207
rect 104 7 120 202
rect 109 2 114 7
rect 119 2 120 7
rect 104 0 120 2
rect 280 307 296 310
rect 285 302 290 307
rect 295 302 296 307
rect 280 107 296 302
rect 285 102 290 107
rect 295 102 296 107
rect 280 0 296 102
use INVX1  INVX1_1
timestamp 1656334919
transform 1 0 4 0 -1 105
box -2 -3 18 103
use OR2X2  OR2X2_1
timestamp 1656334919
transform 1 0 20 0 -1 105
box -2 -3 34 103
use AND2X2  AND2X2_7
timestamp 1656334919
transform -1 0 84 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1656334919
transform -1 0 116 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1656334919
transform 1 0 4 0 1 105
box -2 -3 98 103
use FILL  FILL_1_0_0
timestamp 1656334919
transform 1 0 100 0 1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_2
timestamp 1656334919
transform 1 0 132 0 1 105
box -2 -3 26 103
use INVX1  INVX1_3
timestamp 1656334919
transform 1 0 116 0 1 105
box -2 -3 18 103
use FILL  FILL_1_0_1
timestamp 1656334919
transform 1 0 108 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_5
timestamp 1656334919
transform 1 0 132 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_0_1
timestamp 1656334919
transform 1 0 124 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_0
timestamp 1656334919
transform 1 0 116 0 -1 105
box -2 -3 10 103
use AND2X2  AND2X2_1
timestamp 1656334919
transform -1 0 204 0 1 105
box -2 -3 34 103
use INVX1  INVX1_2
timestamp 1656334919
transform 1 0 156 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_1
timestamp 1656334919
transform -1 0 196 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1656334919
transform 1 0 204 0 1 105
box -2 -3 34 103
use AND2X2  AND2X2_2
timestamp 1656334919
transform -1 0 228 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_2
timestamp 1656334919
transform -1 0 260 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1656334919
transform 1 0 260 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_1_0
timestamp 1656334919
transform 1 0 292 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1656334919
transform 1 0 300 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_1
timestamp 1656334919
transform 1 0 236 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1656334919
transform 1 0 260 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1656334919
transform 1 0 292 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1656334919
transform 1 0 300 0 1 105
box -2 -3 10 103
use AND2X2  AND2X2_4
timestamp 1656334919
transform 1 0 308 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_1
timestamp 1656334919
transform 1 0 340 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1656334919
transform -1 0 388 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1656334919
transform 1 0 388 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1656334919
transform 1 0 308 0 1 105
box -2 -3 98 103
use FILL  FILL_2_1
timestamp 1656334919
transform 1 0 404 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1
timestamp 1656334919
transform -1 0 420 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1656334919
transform 1 0 412 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1656334919
transform 1 0 4 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1656334919
transform -1 0 108 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1656334919
transform -1 0 116 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_6
timestamp 1656334919
transform -1 0 148 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1656334919
transform -1 0 180 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_4
timestamp 1656334919
transform 1 0 180 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_3
timestamp 1656334919
transform -1 0 244 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_3
timestamp 1656334919
transform 1 0 244 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1656334919
transform 1 0 276 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1656334919
transform 1 0 284 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_5
timestamp 1656334919
transform 1 0 292 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1656334919
transform 1 0 324 0 -1 305
box -2 -3 98 103
<< labels >>
flabel metal6 s 104 0 120 8 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 280 0 296 8 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 restart
port 2 nsew
flabel metal3 s -26 68 -22 72 7 FreeSans 24 270 0 0 enable
port 3 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 clk
port 4 nsew
flabel metal3 s 446 48 450 52 3 FreeSans 24 270 0 0 timeout
port 5 nsew
<< end >>
