VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Watchdog
  CLASS BLOCK ;
  FOREIGN Watchdog ;
  ORIGIN 2.600 0.000 ;
  SIZE 47.600 BY 31.000 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 1.400 20.800 1.800 25.000 ;
        RECT 4.200 20.800 4.600 23.100 ;
        RECT 5.800 20.800 6.200 23.100 ;
        RECT 8.600 20.800 9.000 25.100 ;
        RECT 12.600 20.800 13.000 24.900 ;
        RECT 14.200 20.800 14.600 23.100 ;
        RECT 16.100 20.800 16.500 25.100 ;
        RECT 19.000 20.800 19.400 24.500 ;
        RECT 23.000 20.800 23.400 24.500 ;
        RECT 25.900 20.800 26.300 25.100 ;
        RECT 29.400 20.800 29.800 23.100 ;
        RECT 31.000 20.800 31.400 24.900 ;
        RECT 33.400 20.800 33.800 25.000 ;
        RECT 36.200 20.800 36.600 23.100 ;
        RECT 37.800 20.800 38.200 23.100 ;
        RECT 40.600 20.800 41.000 25.100 ;
        RECT 0.200 20.200 42.200 20.800 ;
        RECT 1.400 16.000 1.800 20.200 ;
        RECT 4.200 17.900 4.600 20.200 ;
        RECT 5.800 17.900 6.200 20.200 ;
        RECT 8.600 15.900 9.000 20.200 ;
        RECT 11.800 17.900 12.200 20.200 ;
        RECT 13.400 15.900 13.800 20.200 ;
        RECT 15.800 17.900 16.200 20.200 ;
        RECT 18.200 16.100 18.600 20.200 ;
        RECT 19.800 17.900 20.200 20.200 ;
        RECT 20.600 17.900 21.000 20.200 ;
        RECT 22.200 18.100 22.600 20.200 ;
        RECT 23.800 17.900 24.200 20.200 ;
        RECT 25.400 17.900 25.800 20.200 ;
        RECT 26.200 17.900 26.600 20.200 ;
        RECT 27.800 16.100 28.200 20.200 ;
        RECT 31.800 16.000 32.200 20.200 ;
        RECT 34.600 17.900 35.000 20.200 ;
        RECT 36.200 17.900 36.600 20.200 ;
        RECT 39.000 15.900 39.400 20.200 ;
        RECT 0.600 0.800 1.000 3.100 ;
        RECT 3.500 0.800 3.900 5.100 ;
        RECT 6.200 0.800 6.600 4.900 ;
        RECT 7.800 0.800 8.200 3.100 ;
        RECT 9.700 0.800 10.100 5.100 ;
        RECT 14.200 0.800 14.600 4.500 ;
        RECT 18.200 0.800 18.600 4.500 ;
        RECT 20.600 0.800 21.000 4.900 ;
        RECT 22.200 0.800 22.600 3.100 ;
        RECT 24.600 0.800 25.000 4.500 ;
        RECT 27.500 0.800 27.900 5.100 ;
        RECT 31.000 0.800 31.400 3.100 ;
        RECT 32.600 0.800 33.000 4.900 ;
        RECT 34.200 0.800 34.600 5.100 ;
        RECT 36.600 0.800 37.000 3.100 ;
        RECT 38.200 0.800 38.600 3.100 ;
        RECT 39.800 0.800 40.200 4.500 ;
        RECT 0.200 0.200 42.200 0.800 ;
      LAYER via1 ;
        RECT 10.600 20.300 11.000 20.700 ;
        RECT 11.300 20.300 11.700 20.700 ;
        RECT 10.600 0.300 11.000 0.700 ;
        RECT 11.300 0.300 11.700 0.700 ;
      LAYER metal2 ;
        RECT 10.400 20.300 12.000 20.700 ;
        RECT 10.400 0.300 12.000 0.700 ;
      LAYER via2 ;
        RECT 10.600 20.300 11.000 20.700 ;
        RECT 11.300 20.300 11.700 20.700 ;
        RECT 10.600 0.300 11.000 0.700 ;
        RECT 11.300 0.300 11.700 0.700 ;
      LAYER metal3 ;
        RECT 10.400 20.300 12.000 20.700 ;
        RECT 10.400 0.300 12.000 0.700 ;
      LAYER via3 ;
        RECT 10.600 20.300 11.000 20.700 ;
        RECT 11.400 20.300 11.800 20.700 ;
        RECT 10.600 0.300 11.000 0.700 ;
        RECT 11.400 0.300 11.800 0.700 ;
      LAYER metal4 ;
        RECT 10.400 20.300 12.000 20.700 ;
        RECT 10.400 0.300 12.000 0.700 ;
      LAYER via4 ;
        RECT 10.600 20.300 11.000 20.700 ;
        RECT 11.300 20.300 11.700 20.700 ;
        RECT 10.600 0.300 11.000 0.700 ;
        RECT 11.300 0.300 11.700 0.700 ;
      LAYER metal5 ;
        RECT 10.400 20.200 12.000 20.700 ;
        RECT 10.400 0.200 12.000 0.700 ;
      LAYER via5 ;
        RECT 11.400 20.200 11.900 20.700 ;
        RECT 11.400 0.200 11.900 0.700 ;
      LAYER metal6 ;
        RECT 10.400 0.000 12.000 31.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 30.200 42.200 30.800 ;
        RECT 1.400 27.900 1.800 30.200 ;
        RECT 4.100 28.900 4.600 30.200 ;
        RECT 5.800 28.900 6.200 30.200 ;
        RECT 8.600 28.000 9.000 30.200 ;
        RECT 12.900 28.000 13.300 30.200 ;
        RECT 15.800 28.100 16.200 30.200 ;
        RECT 17.400 28.900 17.800 30.200 ;
        RECT 18.500 27.900 18.900 30.200 ;
        RECT 20.600 28.900 21.000 30.200 ;
        RECT 21.400 28.900 21.800 30.200 ;
        RECT 23.500 27.900 23.900 30.200 ;
        RECT 24.600 28.900 25.000 30.200 ;
        RECT 26.200 28.100 26.600 30.200 ;
        RECT 30.700 28.000 31.100 30.200 ;
        RECT 33.400 27.900 33.800 30.200 ;
        RECT 36.100 28.900 36.600 30.200 ;
        RECT 37.800 28.900 38.200 30.200 ;
        RECT 40.600 28.000 41.000 30.200 ;
        RECT 1.400 10.800 1.800 13.100 ;
        RECT 4.100 10.800 4.600 12.100 ;
        RECT 5.800 10.800 6.200 12.100 ;
        RECT 8.600 10.800 9.000 13.000 ;
        RECT 11.800 10.800 12.200 12.100 ;
        RECT 13.400 10.800 13.800 12.100 ;
        RECT 15.000 10.800 15.400 12.100 ;
        RECT 15.800 10.800 16.200 12.100 ;
        RECT 18.500 10.800 18.900 13.000 ;
        RECT 20.600 10.800 21.000 14.100 ;
        RECT 23.800 10.800 24.200 13.100 ;
        RECT 27.500 10.800 27.900 13.000 ;
        RECT 31.800 10.800 32.200 13.100 ;
        RECT 34.500 10.800 35.000 12.100 ;
        RECT 36.200 10.800 36.600 12.100 ;
        RECT 39.000 10.800 39.400 13.000 ;
        RECT 0.200 10.200 42.200 10.800 ;
        RECT 0.600 8.900 1.000 10.200 ;
        RECT 2.200 8.900 2.600 10.200 ;
        RECT 3.800 8.100 4.200 10.200 ;
        RECT 6.500 8.000 6.900 10.200 ;
        RECT 9.400 8.100 9.800 10.200 ;
        RECT 11.000 8.900 11.400 10.200 ;
        RECT 13.700 7.900 14.100 10.200 ;
        RECT 15.800 8.900 16.200 10.200 ;
        RECT 16.600 8.900 17.000 10.200 ;
        RECT 18.700 7.900 19.100 10.200 ;
        RECT 20.900 8.000 21.300 10.200 ;
        RECT 23.000 8.900 23.400 10.200 ;
        RECT 25.100 7.900 25.500 10.200 ;
        RECT 26.200 8.900 26.600 10.200 ;
        RECT 27.800 8.100 28.200 10.200 ;
        RECT 32.300 8.000 32.700 10.200 ;
        RECT 34.200 8.900 34.600 10.200 ;
        RECT 35.800 8.900 36.200 10.200 ;
        RECT 38.200 7.900 38.600 10.200 ;
        RECT 39.800 7.900 40.200 10.200 ;
      LAYER via1 ;
        RECT 28.200 30.300 28.600 30.700 ;
        RECT 28.900 30.300 29.300 30.700 ;
        RECT 28.200 10.300 28.600 10.700 ;
        RECT 28.900 10.300 29.300 10.700 ;
      LAYER metal2 ;
        RECT 28.000 30.300 29.600 30.700 ;
        RECT 28.000 10.300 29.600 10.700 ;
      LAYER via2 ;
        RECT 28.200 30.300 28.600 30.700 ;
        RECT 28.900 30.300 29.300 30.700 ;
        RECT 28.200 10.300 28.600 10.700 ;
        RECT 28.900 10.300 29.300 10.700 ;
      LAYER metal3 ;
        RECT 28.000 30.300 29.600 30.700 ;
        RECT 28.000 10.300 29.600 10.700 ;
      LAYER via3 ;
        RECT 28.200 30.300 28.600 30.700 ;
        RECT 29.000 30.300 29.400 30.700 ;
        RECT 28.200 10.300 28.600 10.700 ;
        RECT 29.000 10.300 29.400 10.700 ;
      LAYER metal4 ;
        RECT 28.000 30.300 29.600 30.700 ;
        RECT 28.000 10.300 29.600 10.700 ;
      LAYER via4 ;
        RECT 28.200 30.300 28.600 30.700 ;
        RECT 28.900 30.300 29.300 30.700 ;
        RECT 28.200 10.300 28.600 10.700 ;
        RECT 28.900 10.300 29.300 10.700 ;
      LAYER metal5 ;
        RECT 28.000 30.200 29.600 30.700 ;
        RECT 28.000 10.200 29.600 10.700 ;
      LAYER via5 ;
        RECT 29.000 30.200 29.500 30.700 ;
        RECT 29.000 10.200 29.500 10.700 ;
      LAYER metal6 ;
        RECT 28.000 0.000 29.600 31.000 ;
    END
  END gnd
  PIN restart
    PORT
      LAYER metal1 ;
        RECT 3.000 6.800 3.500 7.200 ;
        RECT 3.200 6.400 3.600 6.800 ;
      LAYER metal2 ;
        RECT 3.000 6.800 3.400 7.200 ;
        RECT 3.000 5.200 3.300 6.800 ;
        RECT 3.000 4.800 3.400 5.200 ;
      LAYER metal3 ;
        RECT -2.600 5.100 -2.200 5.200 ;
        RECT 3.000 5.100 3.400 5.200 ;
        RECT -2.600 4.800 3.400 5.100 ;
    END
  END restart
  PIN enable
    PORT
      LAYER metal1 ;
        RECT 0.600 7.800 1.000 8.600 ;
      LAYER metal2 ;
        RECT 0.600 7.800 1.000 8.200 ;
        RECT 0.600 7.200 0.900 7.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
      LAYER metal3 ;
        RECT -2.600 7.100 -2.200 7.200 ;
        RECT 0.600 7.100 1.000 7.200 ;
        RECT -2.600 6.800 1.000 7.100 ;
    END
  END enable
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 3.000 28.200 3.400 28.600 ;
        RECT 35.000 28.200 35.400 28.600 ;
        RECT 1.000 27.100 1.800 27.200 ;
        RECT 3.100 27.100 3.400 28.200 ;
        RECT 35.100 27.200 35.400 28.200 ;
        RECT 5.900 27.100 6.300 27.200 ;
        RECT 33.000 27.100 33.800 27.200 ;
        RECT 35.000 27.100 35.400 27.200 ;
        RECT 37.900 27.100 38.300 27.200 ;
        RECT 1.000 26.800 6.500 27.100 ;
        RECT 33.000 26.800 38.500 27.100 ;
        RECT 2.500 26.700 2.900 26.800 ;
        RECT 6.200 26.200 6.500 26.800 ;
        RECT 34.500 26.700 34.900 26.800 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 6.200 25.200 6.500 25.800 ;
        RECT 38.200 25.200 38.500 26.800 ;
        RECT 6.200 24.900 7.400 25.200 ;
        RECT 38.200 24.900 39.400 25.200 ;
        RECT 7.100 24.400 7.400 24.900 ;
        RECT 39.100 24.400 39.400 24.900 ;
        RECT 7.100 24.000 7.800 24.400 ;
        RECT 39.100 24.000 39.800 24.400 ;
        RECT 7.100 16.600 7.800 17.000 ;
        RECT 37.500 16.600 38.200 17.000 ;
        RECT 7.100 16.100 7.400 16.600 ;
        RECT 37.500 16.100 37.800 16.600 ;
        RECT 6.200 15.800 7.400 16.100 ;
        RECT 36.600 15.800 37.800 16.100 ;
        RECT 6.200 15.200 6.500 15.800 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 2.500 14.200 2.900 14.300 ;
        RECT 6.200 14.200 6.500 14.800 ;
        RECT 32.900 14.200 33.300 14.300 ;
        RECT 36.600 14.200 36.900 15.800 ;
        RECT 1.000 13.900 6.500 14.200 ;
        RECT 31.400 13.900 36.900 14.200 ;
        RECT 1.000 13.800 1.800 13.900 ;
        RECT 3.100 12.800 3.400 13.900 ;
        RECT 5.900 13.800 6.300 13.900 ;
        RECT 31.400 13.800 32.200 13.900 ;
        RECT 33.500 12.800 33.800 13.900 ;
        RECT 35.000 13.800 35.400 13.900 ;
        RECT 36.300 13.800 36.700 13.900 ;
        RECT 3.000 12.400 3.400 12.800 ;
        RECT 33.400 12.400 33.800 12.800 ;
      LAYER via1 ;
        RECT 35.000 26.800 35.400 27.200 ;
      LAYER metal2 ;
        RECT 35.000 26.800 35.400 27.200 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 6.200 16.200 6.500 25.800 ;
        RECT 6.200 15.800 6.600 16.200 ;
        RECT 6.200 15.200 6.500 15.800 ;
        RECT 35.000 15.200 35.300 26.800 ;
        RECT 6.200 14.800 6.600 15.200 ;
        RECT 35.000 14.800 35.400 15.200 ;
        RECT 35.000 14.200 35.300 14.800 ;
        RECT 35.000 13.800 35.400 14.200 ;
      LAYER metal3 ;
        RECT 6.200 15.800 6.600 16.200 ;
        RECT -2.600 15.100 -2.200 15.200 ;
        RECT 6.200 15.100 6.500 15.800 ;
        RECT 35.000 15.100 35.400 15.200 ;
        RECT -2.600 14.800 35.400 15.100 ;
    END
  END clk
  PIN timeout
    PORT
      LAYER metal1 ;
        RECT 40.600 6.200 41.000 9.900 ;
        RECT 40.700 5.100 41.000 6.200 ;
        RECT 40.600 4.100 41.000 5.100 ;
        RECT 41.400 4.100 41.800 4.200 ;
        RECT 40.600 3.800 41.800 4.100 ;
        RECT 40.600 1.100 41.000 3.800 ;
      LAYER via1 ;
        RECT 41.400 3.800 41.800 4.200 ;
      LAYER metal2 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 41.400 4.200 41.700 4.800 ;
        RECT 41.400 3.800 41.800 4.200 ;
      LAYER metal3 ;
        RECT 41.400 5.100 41.800 5.200 ;
        RECT 44.600 5.100 45.000 5.200 ;
        RECT 41.400 4.800 45.000 5.100 ;
    END
  END timeout
  OBS
      LAYER metal1 ;
        RECT 0.600 27.500 1.000 29.900 ;
        RECT 2.800 29.200 3.200 29.900 ;
        RECT 2.200 28.900 3.200 29.200 ;
        RECT 5.000 28.900 5.400 29.900 ;
        RECT 7.100 29.200 7.700 29.900 ;
        RECT 7.000 28.900 7.700 29.200 ;
        RECT 2.200 28.500 2.600 28.900 ;
        RECT 5.000 28.600 5.300 28.900 ;
        RECT 3.900 28.300 5.300 28.600 ;
        RECT 7.000 28.500 7.400 28.900 ;
        RECT 3.900 28.200 4.300 28.300 ;
        RECT 7.900 27.700 8.300 27.800 ;
        RECT 9.400 27.700 9.800 29.900 ;
        RECT 12.100 28.400 12.500 29.900 ;
        RECT 7.900 27.400 9.800 27.700 ;
        RECT 7.000 26.400 7.400 26.500 ;
        RECT 1.700 26.200 2.100 26.300 ;
        RECT 1.700 25.900 4.200 26.200 ;
        RECT 7.000 26.100 8.900 26.400 ;
        RECT 8.500 26.000 8.900 26.100 ;
        RECT 3.800 25.800 4.200 25.900 ;
        RECT 7.700 25.700 8.100 25.800 ;
        RECT 9.400 25.700 9.800 27.400 ;
        RECT 11.800 27.900 12.500 28.400 ;
        RECT 14.200 27.900 14.600 29.900 ;
        RECT 15.000 27.900 15.400 29.900 ;
        RECT 16.600 28.900 17.000 29.900 ;
        RECT 11.800 26.200 12.100 27.900 ;
        RECT 14.200 27.800 14.500 27.900 ;
        RECT 13.600 27.600 14.500 27.800 ;
        RECT 12.400 27.500 14.500 27.600 ;
        RECT 12.400 27.300 13.900 27.500 ;
        RECT 12.400 27.200 12.800 27.300 ;
        RECT 11.000 26.100 11.400 26.200 ;
        RECT 11.800 26.100 12.200 26.200 ;
        RECT 11.000 25.800 12.200 26.100 ;
        RECT 0.600 25.500 3.400 25.600 ;
        RECT 0.600 25.400 3.500 25.500 ;
        RECT 7.700 25.400 9.800 25.700 ;
        RECT 0.600 25.300 5.500 25.400 ;
        RECT 0.600 21.100 1.000 25.300 ;
        RECT 3.100 25.100 5.500 25.300 ;
        RECT 2.200 24.500 4.900 24.800 ;
        RECT 2.200 24.400 2.600 24.500 ;
        RECT 4.500 24.400 4.900 24.500 ;
        RECT 5.200 24.500 5.500 25.100 ;
        RECT 5.900 24.500 6.300 24.600 ;
        RECT 5.200 24.200 6.300 24.500 ;
        RECT 3.900 23.700 4.300 23.800 ;
        RECT 5.300 23.700 5.700 23.800 ;
        RECT 2.200 23.100 2.600 23.500 ;
        RECT 3.900 23.400 5.700 23.700 ;
        RECT 5.000 23.100 5.300 23.400 ;
        RECT 7.000 23.100 7.400 23.500 ;
        RECT 2.200 22.800 3.200 23.100 ;
        RECT 2.800 21.100 3.200 22.800 ;
        RECT 5.000 21.100 5.400 23.100 ;
        RECT 7.100 21.100 7.700 23.100 ;
        RECT 9.400 21.100 9.800 25.400 ;
        RECT 11.800 25.100 12.100 25.800 ;
        RECT 12.500 25.500 12.800 27.200 ;
        RECT 14.200 27.100 14.600 27.200 ;
        RECT 15.000 27.100 15.300 27.900 ;
        RECT 16.600 27.800 16.900 28.900 ;
        RECT 17.400 27.800 17.800 28.600 ;
        RECT 19.800 27.800 20.200 29.900 ;
        RECT 20.500 28.200 20.900 28.600 ;
        RECT 21.500 28.200 21.900 28.600 ;
        RECT 20.600 28.100 21.000 28.200 ;
        RECT 21.400 28.100 21.800 28.200 ;
        RECT 20.600 27.800 21.800 28.100 ;
        RECT 22.200 27.900 22.600 29.900 ;
        RECT 25.400 28.900 25.800 29.900 ;
        RECT 13.200 26.600 13.800 27.000 ;
        RECT 14.200 26.800 15.300 27.100 ;
        RECT 13.400 26.200 13.700 26.600 ;
        RECT 14.200 26.400 14.600 26.800 ;
        RECT 15.000 26.200 15.300 26.800 ;
        RECT 15.700 27.500 16.900 27.800 ;
        RECT 13.400 25.800 13.800 26.200 ;
        RECT 15.000 25.800 15.400 26.200 ;
        RECT 15.700 26.000 16.000 27.500 ;
        RECT 16.500 27.100 17.000 27.200 ;
        RECT 19.000 27.100 19.400 27.200 ;
        RECT 16.500 26.800 19.400 27.100 ;
        RECT 16.400 26.400 16.800 26.800 ;
        RECT 19.000 26.400 19.400 26.800 ;
        RECT 18.200 26.100 18.600 26.200 ;
        RECT 19.800 26.100 20.100 27.800 ;
        RECT 22.300 26.200 22.600 27.900 ;
        RECT 24.600 27.800 25.000 28.600 ;
        RECT 25.500 27.800 25.800 28.900 ;
        RECT 27.000 27.900 27.400 29.900 ;
        RECT 29.400 27.900 29.800 29.900 ;
        RECT 31.500 28.400 31.900 29.900 ;
        RECT 31.500 27.900 32.200 28.400 ;
        RECT 25.500 27.500 26.700 27.800 ;
        RECT 23.000 27.100 23.400 27.200 ;
        RECT 25.400 27.100 25.900 27.200 ;
        RECT 23.000 26.800 25.900 27.100 ;
        RECT 23.000 26.400 23.400 26.800 ;
        RECT 25.600 26.400 26.000 26.800 ;
        RECT 20.600 26.100 21.000 26.200 ;
        RECT 12.500 25.200 13.700 25.500 ;
        RECT 11.800 21.100 12.200 25.100 ;
        RECT 13.400 23.100 13.700 25.200 ;
        RECT 15.000 25.100 15.300 25.800 ;
        RECT 15.700 25.700 16.100 26.000 ;
        RECT 18.200 25.800 19.000 26.100 ;
        RECT 19.800 25.800 21.000 26.100 ;
        RECT 21.400 26.100 21.800 26.200 ;
        RECT 22.200 26.100 22.600 26.200 ;
        RECT 23.800 26.100 24.200 26.200 ;
        RECT 21.400 25.800 22.600 26.100 ;
        RECT 23.400 25.800 24.200 26.100 ;
        RECT 26.400 26.000 26.700 27.500 ;
        RECT 27.100 27.100 27.400 27.900 ;
        RECT 29.500 27.800 29.800 27.900 ;
        RECT 29.500 27.600 30.400 27.800 ;
        RECT 29.500 27.500 31.600 27.600 ;
        RECT 30.100 27.300 31.600 27.500 ;
        RECT 31.200 27.200 31.600 27.300 ;
        RECT 29.400 27.100 29.800 27.200 ;
        RECT 27.000 26.800 29.800 27.100 ;
        RECT 30.400 26.900 30.800 27.000 ;
        RECT 27.100 26.200 27.400 26.800 ;
        RECT 29.400 26.400 29.800 26.800 ;
        RECT 30.300 26.600 30.800 26.900 ;
        RECT 30.300 26.200 30.600 26.600 ;
        RECT 15.700 25.600 17.800 25.700 ;
        RECT 18.600 25.600 19.000 25.800 ;
        RECT 15.800 25.400 17.800 25.600 ;
        RECT 15.000 24.800 15.700 25.100 ;
        RECT 13.400 21.100 13.800 23.100 ;
        RECT 15.300 21.100 15.700 24.800 ;
        RECT 17.400 21.100 17.800 25.400 ;
        RECT 20.600 25.100 20.900 25.800 ;
        RECT 21.500 25.100 21.800 25.800 ;
        RECT 23.400 25.600 23.800 25.800 ;
        RECT 26.300 25.700 26.700 26.000 ;
        RECT 27.000 25.800 27.400 26.200 ;
        RECT 30.200 25.800 30.600 26.200 ;
        RECT 24.600 25.600 26.700 25.700 ;
        RECT 24.600 25.400 26.600 25.600 ;
        RECT 18.200 24.800 20.200 25.100 ;
        RECT 18.200 21.100 18.600 24.800 ;
        RECT 19.800 21.100 20.200 24.800 ;
        RECT 20.600 21.100 21.000 25.100 ;
        RECT 21.400 21.100 21.800 25.100 ;
        RECT 22.200 24.800 24.200 25.100 ;
        RECT 22.200 21.100 22.600 24.800 ;
        RECT 23.800 21.100 24.200 24.800 ;
        RECT 24.600 21.100 25.000 25.400 ;
        RECT 27.100 25.100 27.400 25.800 ;
        RECT 31.200 25.500 31.500 27.200 ;
        RECT 31.900 26.200 32.200 27.900 ;
        RECT 32.600 27.500 33.000 29.900 ;
        RECT 34.800 29.200 35.200 29.900 ;
        RECT 34.200 28.900 35.200 29.200 ;
        RECT 37.000 28.900 37.400 29.900 ;
        RECT 39.100 29.200 39.700 29.900 ;
        RECT 39.000 28.900 39.700 29.200 ;
        RECT 34.200 28.500 34.600 28.900 ;
        RECT 37.000 28.600 37.300 28.900 ;
        RECT 35.900 28.300 37.300 28.600 ;
        RECT 39.000 28.500 39.400 28.900 ;
        RECT 35.900 28.200 36.300 28.300 ;
        RECT 39.900 27.700 40.300 27.800 ;
        RECT 41.400 27.700 41.800 29.900 ;
        RECT 39.900 27.400 41.800 27.700 ;
        RECT 39.000 26.400 39.400 26.500 ;
        RECT 31.800 25.800 32.200 26.200 ;
        RECT 33.700 26.200 34.100 26.300 ;
        RECT 33.700 25.900 36.200 26.200 ;
        RECT 39.000 26.100 40.900 26.400 ;
        RECT 40.500 26.000 40.900 26.100 ;
        RECT 35.800 25.800 36.200 25.900 ;
        RECT 26.700 24.800 27.400 25.100 ;
        RECT 30.300 25.200 31.500 25.500 ;
        RECT 26.700 21.100 27.100 24.800 ;
        RECT 30.300 23.100 30.600 25.200 ;
        RECT 31.900 25.100 32.200 25.800 ;
        RECT 39.700 25.700 40.100 25.800 ;
        RECT 41.400 25.700 41.800 27.400 ;
        RECT 30.200 21.100 30.600 23.100 ;
        RECT 31.800 21.100 32.200 25.100 ;
        RECT 32.600 25.500 35.400 25.600 ;
        RECT 32.600 25.400 35.500 25.500 ;
        RECT 39.700 25.400 41.800 25.700 ;
        RECT 32.600 25.300 37.500 25.400 ;
        RECT 32.600 21.100 33.000 25.300 ;
        RECT 35.100 25.100 37.500 25.300 ;
        RECT 34.200 24.500 36.900 24.800 ;
        RECT 34.200 24.400 34.600 24.500 ;
        RECT 36.500 24.400 36.900 24.500 ;
        RECT 37.200 24.500 37.500 25.100 ;
        RECT 37.900 24.500 38.300 24.600 ;
        RECT 37.200 24.200 38.300 24.500 ;
        RECT 35.900 23.700 36.300 23.800 ;
        RECT 37.300 23.700 37.700 23.800 ;
        RECT 34.200 23.100 34.600 23.500 ;
        RECT 35.900 23.400 37.700 23.700 ;
        RECT 37.000 23.100 37.300 23.400 ;
        RECT 39.000 23.100 39.400 23.500 ;
        RECT 34.200 22.800 35.200 23.100 ;
        RECT 34.800 21.100 35.200 22.800 ;
        RECT 37.000 21.100 37.400 23.100 ;
        RECT 39.100 21.100 39.700 23.100 ;
        RECT 41.400 21.100 41.800 25.400 ;
        RECT 0.600 15.700 1.000 19.900 ;
        RECT 2.800 18.200 3.200 19.900 ;
        RECT 2.200 17.900 3.200 18.200 ;
        RECT 5.000 17.900 5.400 19.900 ;
        RECT 7.100 17.900 7.700 19.900 ;
        RECT 2.200 17.500 2.600 17.900 ;
        RECT 5.000 17.600 5.300 17.900 ;
        RECT 3.900 17.300 5.700 17.600 ;
        RECT 7.000 17.500 7.400 17.900 ;
        RECT 3.900 17.200 4.300 17.300 ;
        RECT 5.300 17.200 5.700 17.300 ;
        RECT 2.200 16.500 2.600 16.600 ;
        RECT 4.500 16.500 4.900 16.600 ;
        RECT 2.200 16.200 4.900 16.500 ;
        RECT 5.200 16.500 6.300 16.800 ;
        RECT 5.200 15.900 5.500 16.500 ;
        RECT 5.900 16.400 6.300 16.500 ;
        RECT 3.100 15.700 5.500 15.900 ;
        RECT 0.600 15.600 5.500 15.700 ;
        RECT 9.400 15.600 9.800 19.900 ;
        RECT 0.600 15.500 3.500 15.600 ;
        RECT 0.600 15.400 3.400 15.500 ;
        RECT 7.700 15.300 9.800 15.600 ;
        RECT 7.700 15.200 8.100 15.300 ;
        RECT 3.800 15.100 4.200 15.200 ;
        RECT 5.400 15.100 5.800 15.200 ;
        RECT 1.700 14.800 5.800 15.100 ;
        RECT 8.500 14.900 8.900 15.000 ;
        RECT 1.700 14.700 2.100 14.800 ;
        RECT 7.000 14.600 8.900 14.900 ;
        RECT 7.000 14.500 7.400 14.600 ;
        RECT 9.400 13.600 9.800 15.300 ;
        RECT 0.600 11.100 1.000 13.500 ;
        RECT 7.900 13.300 9.800 13.600 ;
        RECT 7.900 13.200 8.300 13.300 ;
        RECT 3.900 12.700 4.300 12.800 ;
        RECT 2.200 12.100 2.600 12.500 ;
        RECT 3.900 12.400 5.300 12.700 ;
        RECT 5.000 12.100 5.300 12.400 ;
        RECT 7.000 12.100 7.400 12.500 ;
        RECT 9.400 12.100 9.800 13.300 ;
        RECT 11.800 12.400 12.200 13.200 ;
        RECT 12.600 13.100 13.000 19.900 ;
        RECT 14.700 16.300 15.100 19.900 ;
        RECT 14.200 15.900 15.100 16.300 ;
        RECT 14.300 14.200 14.600 15.900 ;
        RECT 15.000 15.100 15.400 15.600 ;
        RECT 15.800 15.100 16.200 15.200 ;
        RECT 15.000 14.800 16.200 15.100 ;
        RECT 13.400 14.100 13.800 14.200 ;
        RECT 14.200 14.100 14.600 14.200 ;
        RECT 13.400 13.800 14.600 14.100 ;
        RECT 13.400 13.100 13.800 13.200 ;
        RECT 12.600 12.800 13.800 13.100 ;
        RECT 10.200 12.100 10.600 12.200 ;
        RECT 2.200 11.800 3.200 12.100 ;
        RECT 2.800 11.100 3.200 11.800 ;
        RECT 5.000 11.100 5.400 12.100 ;
        RECT 7.000 11.800 7.700 12.100 ;
        RECT 7.100 11.100 7.700 11.800 ;
        RECT 9.400 11.800 10.600 12.100 ;
        RECT 9.400 11.100 9.800 11.800 ;
        RECT 12.600 11.100 13.000 12.800 ;
        RECT 13.400 12.400 13.800 12.800 ;
        RECT 14.300 12.100 14.600 13.800 ;
        RECT 15.800 12.400 16.200 13.200 ;
        RECT 14.200 11.100 14.600 12.100 ;
        RECT 16.600 11.100 17.000 19.900 ;
        RECT 17.400 15.900 17.800 19.900 ;
        RECT 19.000 17.900 19.400 19.900 ;
        RECT 21.400 17.900 21.800 19.900 ;
        RECT 17.400 15.200 17.700 15.900 ;
        RECT 19.000 15.800 19.300 17.900 ;
        RECT 21.500 17.800 21.800 17.900 ;
        RECT 23.000 17.900 23.400 19.900 ;
        RECT 23.000 17.800 23.300 17.900 ;
        RECT 21.500 17.500 23.300 17.800 ;
        RECT 22.200 16.400 22.600 17.200 ;
        RECT 23.000 16.200 23.300 17.500 ;
        RECT 18.100 15.500 19.300 15.800 ;
        RECT 17.400 14.800 17.800 15.200 ;
        RECT 17.400 13.100 17.700 14.800 ;
        RECT 18.100 13.800 18.400 15.500 ;
        RECT 20.600 15.400 21.000 16.200 ;
        RECT 23.000 15.800 23.400 16.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 21.400 14.800 22.200 15.200 ;
        RECT 19.000 14.400 19.300 14.800 ;
        RECT 18.800 14.100 19.300 14.400 ;
        RECT 18.800 14.000 19.200 14.100 ;
        RECT 19.800 13.800 20.200 14.600 ;
        RECT 23.000 14.200 23.300 15.800 ;
        RECT 22.500 14.100 23.300 14.200 ;
        RECT 22.400 13.900 23.300 14.100 ;
        RECT 18.000 13.700 18.400 13.800 ;
        RECT 18.000 13.500 19.500 13.700 ;
        RECT 18.000 13.400 20.100 13.500 ;
        RECT 19.200 13.200 20.100 13.400 ;
        RECT 22.400 13.200 22.800 13.900 ;
        RECT 23.800 13.400 24.200 14.200 ;
        RECT 19.800 13.100 20.100 13.200 ;
        RECT 17.400 12.600 18.100 13.100 ;
        RECT 17.700 12.200 18.100 12.600 ;
        RECT 17.400 11.800 18.100 12.200 ;
        RECT 17.700 11.100 18.100 11.800 ;
        RECT 19.800 11.100 20.200 13.100 ;
        RECT 22.200 12.800 22.800 13.200 ;
        RECT 24.600 13.100 25.000 19.900 ;
        RECT 27.000 17.900 27.400 19.900 ;
        RECT 25.400 15.800 25.800 16.600 ;
        RECT 27.100 15.800 27.400 17.900 ;
        RECT 28.600 19.100 29.000 19.900 ;
        RECT 29.400 19.100 29.800 19.200 ;
        RECT 28.600 18.800 29.800 19.100 ;
        RECT 28.600 15.900 29.000 18.800 ;
        RECT 27.100 15.500 28.300 15.800 ;
        RECT 27.000 14.800 27.400 15.200 ;
        RECT 26.200 13.800 26.600 14.600 ;
        RECT 27.100 14.400 27.400 14.800 ;
        RECT 27.100 14.100 27.600 14.400 ;
        RECT 27.200 14.000 27.600 14.100 ;
        RECT 28.000 13.800 28.300 15.500 ;
        RECT 28.700 15.200 29.000 15.900 ;
        RECT 31.000 15.700 31.400 19.900 ;
        RECT 33.200 18.200 33.600 19.900 ;
        RECT 32.600 17.900 33.600 18.200 ;
        RECT 35.400 17.900 35.800 19.900 ;
        RECT 37.500 17.900 38.100 19.900 ;
        RECT 32.600 17.500 33.000 17.900 ;
        RECT 35.400 17.600 35.700 17.900 ;
        RECT 34.300 17.300 36.100 17.600 ;
        RECT 37.400 17.500 37.800 17.900 ;
        RECT 34.300 17.200 34.700 17.300 ;
        RECT 35.700 17.200 36.100 17.300 ;
        RECT 32.600 16.500 33.000 16.600 ;
        RECT 34.900 16.500 35.300 16.600 ;
        RECT 32.600 16.200 35.300 16.500 ;
        RECT 35.600 16.500 36.700 16.800 ;
        RECT 35.600 15.900 35.900 16.500 ;
        RECT 36.300 16.400 36.700 16.500 ;
        RECT 33.500 15.700 35.900 15.900 ;
        RECT 31.000 15.600 35.900 15.700 ;
        RECT 39.800 15.600 40.200 19.900 ;
        RECT 31.000 15.500 33.900 15.600 ;
        RECT 31.000 15.400 33.800 15.500 ;
        RECT 38.100 15.300 40.200 15.600 ;
        RECT 38.100 15.200 38.500 15.300 ;
        RECT 28.600 14.800 29.000 15.200 ;
        RECT 34.200 15.100 34.600 15.200 ;
        RECT 28.000 13.700 28.400 13.800 ;
        RECT 26.900 13.500 28.400 13.700 ;
        RECT 26.300 13.400 28.400 13.500 ;
        RECT 26.300 13.200 27.200 13.400 ;
        RECT 26.300 13.100 26.600 13.200 ;
        RECT 28.700 13.100 29.000 14.800 ;
        RECT 32.100 14.800 34.600 15.100 ;
        RECT 38.900 14.900 39.300 15.000 ;
        RECT 32.100 14.700 32.500 14.800 ;
        RECT 33.400 14.700 33.800 14.800 ;
        RECT 37.400 14.600 39.300 14.900 ;
        RECT 37.400 14.500 37.800 14.600 ;
        RECT 39.800 13.600 40.200 15.300 ;
        RECT 24.600 12.800 25.500 13.100 ;
        RECT 22.400 11.100 22.800 12.800 ;
        RECT 25.100 12.200 25.500 12.800 ;
        RECT 24.600 11.800 25.500 12.200 ;
        RECT 25.100 11.100 25.500 11.800 ;
        RECT 26.200 11.100 26.600 13.100 ;
        RECT 28.300 12.600 29.000 13.100 ;
        RECT 28.300 11.100 28.700 12.600 ;
        RECT 31.000 11.100 31.400 13.500 ;
        RECT 38.300 13.300 40.200 13.600 ;
        RECT 38.300 13.200 38.700 13.300 ;
        RECT 34.300 12.700 34.700 12.800 ;
        RECT 32.600 12.100 33.000 12.500 ;
        RECT 34.300 12.400 35.700 12.700 ;
        RECT 35.400 12.100 35.700 12.400 ;
        RECT 37.400 12.100 37.800 12.500 ;
        RECT 32.600 11.800 33.600 12.100 ;
        RECT 33.200 11.100 33.600 11.800 ;
        RECT 35.400 11.100 35.800 12.100 ;
        RECT 37.400 11.800 38.100 12.100 ;
        RECT 37.500 11.100 38.100 11.800 ;
        RECT 39.800 11.100 40.200 13.300 ;
        RECT 1.400 8.100 1.800 9.900 ;
        RECT 3.000 8.900 3.400 9.900 ;
        RECT 2.200 8.100 2.600 8.600 ;
        RECT 1.400 7.800 2.600 8.100 ;
        RECT 3.100 7.800 3.400 8.900 ;
        RECT 4.600 7.900 5.000 9.900 ;
        RECT 5.700 9.200 6.100 9.900 ;
        RECT 5.400 8.800 6.100 9.200 ;
        RECT 5.700 8.400 6.100 8.800 ;
        RECT 1.400 7.100 1.800 7.800 ;
        RECT 3.100 7.500 4.300 7.800 ;
        RECT 2.200 7.100 2.600 7.200 ;
        RECT 1.400 6.800 2.600 7.100 ;
        RECT 1.400 1.100 1.800 6.800 ;
        RECT 4.000 6.000 4.300 7.500 ;
        RECT 4.700 6.200 5.000 7.900 ;
        RECT 3.900 5.700 4.300 6.000 ;
        RECT 4.600 5.800 5.000 6.200 ;
        RECT 2.200 5.600 4.300 5.700 ;
        RECT 2.200 5.400 4.200 5.600 ;
        RECT 2.200 1.100 2.600 5.400 ;
        RECT 4.700 5.100 5.000 5.800 ;
        RECT 4.300 4.800 5.000 5.100 ;
        RECT 5.400 7.900 6.100 8.400 ;
        RECT 7.800 7.900 8.200 9.900 ;
        RECT 8.600 7.900 9.000 9.900 ;
        RECT 10.200 8.900 10.600 9.900 ;
        RECT 5.400 6.200 5.700 7.900 ;
        RECT 7.800 7.800 8.100 7.900 ;
        RECT 7.200 7.600 8.100 7.800 ;
        RECT 6.000 7.500 8.100 7.600 ;
        RECT 6.000 7.300 7.500 7.500 ;
        RECT 6.000 7.200 6.400 7.300 ;
        RECT 5.400 5.800 5.800 6.200 ;
        RECT 5.400 5.100 5.700 5.800 ;
        RECT 6.100 5.500 6.400 7.200 ;
        RECT 7.800 7.100 8.200 7.200 ;
        RECT 8.600 7.100 8.900 7.900 ;
        RECT 10.200 7.800 10.500 8.900 ;
        RECT 11.000 8.100 11.400 8.600 ;
        RECT 11.800 8.100 12.200 8.200 ;
        RECT 11.000 7.800 12.200 8.100 ;
        RECT 15.000 7.800 15.400 9.900 ;
        RECT 15.700 8.200 16.100 8.600 ;
        RECT 16.700 8.200 17.100 8.600 ;
        RECT 15.800 7.800 16.200 8.200 ;
        RECT 16.600 7.800 17.000 8.200 ;
        RECT 17.400 7.900 17.800 9.900 ;
        RECT 20.100 8.400 20.500 9.900 ;
        RECT 6.800 6.900 7.200 7.000 ;
        RECT 6.800 6.600 7.300 6.900 ;
        RECT 7.000 6.200 7.300 6.600 ;
        RECT 7.800 6.800 8.900 7.100 ;
        RECT 7.800 6.400 8.200 6.800 ;
        RECT 8.600 6.200 8.900 6.800 ;
        RECT 9.300 7.500 10.500 7.800 ;
        RECT 7.000 5.800 7.400 6.200 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 9.300 6.000 9.600 7.500 ;
        RECT 10.100 7.100 10.600 7.200 ;
        RECT 14.200 7.100 14.600 7.200 ;
        RECT 10.100 6.800 14.600 7.100 ;
        RECT 10.000 6.400 10.400 6.800 ;
        RECT 14.200 6.400 14.600 6.800 ;
        RECT 11.800 6.100 12.200 6.200 ;
        RECT 13.400 6.100 13.800 6.200 ;
        RECT 15.000 6.100 15.300 7.800 ;
        RECT 15.800 6.100 16.200 6.200 ;
        RECT 6.100 5.200 7.300 5.500 ;
        RECT 4.300 1.100 4.700 4.800 ;
        RECT 5.400 1.100 5.800 5.100 ;
        RECT 7.000 3.100 7.300 5.200 ;
        RECT 8.600 5.100 8.900 5.800 ;
        RECT 9.300 5.700 9.700 6.000 ;
        RECT 11.800 5.800 14.200 6.100 ;
        RECT 15.000 5.800 16.200 6.100 ;
        RECT 16.600 6.100 17.000 6.200 ;
        RECT 17.500 6.100 17.800 7.900 ;
        RECT 19.800 7.900 20.500 8.400 ;
        RECT 22.200 7.900 22.600 9.900 ;
        RECT 23.100 8.200 23.500 8.600 ;
        RECT 18.200 7.100 18.600 7.200 ;
        RECT 19.000 7.100 19.400 7.200 ;
        RECT 18.200 6.800 19.400 7.100 ;
        RECT 18.200 6.400 18.600 6.800 ;
        RECT 19.800 6.200 20.100 7.900 ;
        RECT 22.200 7.800 22.500 7.900 ;
        RECT 23.000 7.800 23.400 8.200 ;
        RECT 23.800 7.900 24.200 9.900 ;
        RECT 27.000 8.900 27.400 9.900 ;
        RECT 21.600 7.600 22.500 7.800 ;
        RECT 20.400 7.500 22.500 7.600 ;
        RECT 20.400 7.300 21.900 7.500 ;
        RECT 20.400 7.200 20.800 7.300 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 16.600 5.800 17.800 6.100 ;
        RECT 18.600 5.800 19.400 6.100 ;
        RECT 19.800 5.800 20.200 6.200 ;
        RECT 9.300 5.600 11.400 5.700 ;
        RECT 13.800 5.600 14.200 5.800 ;
        RECT 9.400 5.400 11.400 5.600 ;
        RECT 8.600 4.800 9.300 5.100 ;
        RECT 7.000 1.100 7.400 3.100 ;
        RECT 8.900 1.100 9.300 4.800 ;
        RECT 11.000 1.100 11.400 5.400 ;
        RECT 15.800 5.100 16.100 5.800 ;
        RECT 16.700 5.100 17.000 5.800 ;
        RECT 18.600 5.600 19.000 5.800 ;
        RECT 19.800 5.100 20.100 5.800 ;
        RECT 20.500 5.500 20.800 7.200 ;
        RECT 22.200 7.100 22.600 7.200 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 21.200 6.600 21.800 7.000 ;
        RECT 22.200 6.800 23.400 7.100 ;
        RECT 21.400 6.200 21.700 6.600 ;
        RECT 22.200 6.400 22.600 6.800 ;
        RECT 23.900 6.200 24.200 7.900 ;
        RECT 26.200 7.800 26.600 8.600 ;
        RECT 27.100 7.800 27.400 8.900 ;
        RECT 28.600 7.900 29.000 9.900 ;
        RECT 31.000 7.900 31.400 9.900 ;
        RECT 33.100 9.200 33.500 9.900 ;
        RECT 33.100 8.800 33.800 9.200 ;
        RECT 35.000 8.900 35.400 9.900 ;
        RECT 33.100 8.400 33.500 8.800 ;
        RECT 33.100 7.900 33.800 8.400 ;
        RECT 27.100 7.500 28.300 7.800 ;
        RECT 24.600 7.100 25.000 7.200 ;
        RECT 27.000 7.100 27.500 7.200 ;
        RECT 24.600 6.800 27.500 7.100 ;
        RECT 24.600 6.400 25.000 6.800 ;
        RECT 27.200 6.400 27.600 6.800 ;
        RECT 21.400 5.800 21.800 6.200 ;
        RECT 23.000 6.100 23.400 6.200 ;
        RECT 23.800 6.100 24.200 6.200 ;
        RECT 25.400 6.100 25.800 6.200 ;
        RECT 23.000 5.800 24.200 6.100 ;
        RECT 25.000 5.800 25.800 6.100 ;
        RECT 28.000 6.000 28.300 7.500 ;
        RECT 28.700 7.100 29.000 7.900 ;
        RECT 31.100 7.800 31.400 7.900 ;
        RECT 31.100 7.600 32.000 7.800 ;
        RECT 31.100 7.500 33.200 7.600 ;
        RECT 31.700 7.300 33.200 7.500 ;
        RECT 32.800 7.200 33.200 7.300 ;
        RECT 31.000 7.100 31.400 7.200 ;
        RECT 28.600 6.800 31.400 7.100 ;
        RECT 32.000 6.900 32.400 7.000 ;
        RECT 28.700 6.200 29.000 6.800 ;
        RECT 31.000 6.400 31.400 6.800 ;
        RECT 31.900 6.600 32.400 6.900 ;
        RECT 31.900 6.200 32.200 6.600 ;
        RECT 20.500 5.200 21.700 5.500 ;
        RECT 13.400 4.800 15.400 5.100 ;
        RECT 13.400 1.100 13.800 4.800 ;
        RECT 15.000 1.100 15.400 4.800 ;
        RECT 15.800 1.100 16.200 5.100 ;
        RECT 16.600 1.100 17.000 5.100 ;
        RECT 17.400 4.800 19.400 5.100 ;
        RECT 17.400 1.100 17.800 4.800 ;
        RECT 19.000 1.100 19.400 4.800 ;
        RECT 19.800 1.100 20.200 5.100 ;
        RECT 21.400 3.100 21.700 5.200 ;
        RECT 23.100 5.100 23.400 5.800 ;
        RECT 25.000 5.600 25.400 5.800 ;
        RECT 27.900 5.700 28.300 6.000 ;
        RECT 28.600 5.800 29.000 6.200 ;
        RECT 31.800 5.800 32.200 6.200 ;
        RECT 26.200 5.600 28.300 5.700 ;
        RECT 26.200 5.400 28.200 5.600 ;
        RECT 21.400 1.100 21.800 3.100 ;
        RECT 23.000 1.100 23.400 5.100 ;
        RECT 23.800 4.800 25.800 5.100 ;
        RECT 23.800 1.100 24.200 4.800 ;
        RECT 25.400 1.100 25.800 4.800 ;
        RECT 26.200 1.100 26.600 5.400 ;
        RECT 28.700 5.100 29.000 5.800 ;
        RECT 32.800 5.500 33.100 7.200 ;
        RECT 33.500 6.200 33.800 7.900 ;
        RECT 34.200 7.800 34.600 8.600 ;
        RECT 35.100 7.200 35.400 8.900 ;
        RECT 36.900 8.200 37.300 9.900 ;
        RECT 36.900 7.900 37.800 8.200 ;
        RECT 35.000 6.800 35.400 7.200 ;
        RECT 33.400 5.800 33.800 6.200 ;
        RECT 34.200 6.100 34.600 6.200 ;
        RECT 35.100 6.100 35.400 6.800 ;
        RECT 34.200 5.800 35.400 6.100 ;
        RECT 28.300 4.800 29.000 5.100 ;
        RECT 31.900 5.200 33.100 5.500 ;
        RECT 28.300 1.100 28.700 4.800 ;
        RECT 31.900 3.100 32.200 5.200 ;
        RECT 33.500 5.100 33.800 5.800 ;
        RECT 35.100 5.100 35.400 5.800 ;
        RECT 35.800 6.100 36.200 6.200 ;
        RECT 37.400 6.100 37.800 7.900 ;
        RECT 39.000 7.600 39.400 9.900 ;
        RECT 38.200 6.800 38.600 7.600 ;
        RECT 39.000 7.300 40.100 7.600 ;
        RECT 35.800 5.800 37.800 6.100 ;
        RECT 39.000 5.800 39.400 6.600 ;
        RECT 39.800 5.800 40.100 7.300 ;
        RECT 35.800 5.400 36.200 5.800 ;
        RECT 31.800 1.100 32.200 3.100 ;
        RECT 33.400 1.100 33.800 5.100 ;
        RECT 35.000 4.700 35.900 5.100 ;
        RECT 35.500 1.100 35.900 4.700 ;
        RECT 36.600 4.400 37.000 5.200 ;
        RECT 37.400 1.100 37.800 5.800 ;
        RECT 39.800 5.400 40.400 5.800 ;
        RECT 39.800 5.100 40.100 5.400 ;
        RECT 39.000 4.800 40.100 5.100 ;
        RECT 39.000 1.100 39.400 4.800 ;
      LAYER via1 ;
        RECT 0.600 25.100 1.000 25.500 ;
        RECT 9.400 21.800 9.800 22.200 ;
        RECT 13.400 26.600 13.800 27.000 ;
        RECT 19.000 26.800 19.400 27.200 ;
        RECT 22.200 25.800 22.600 26.200 ;
        RECT 23.800 25.800 24.200 26.200 ;
        RECT 32.600 25.100 33.000 25.500 ;
        RECT 41.400 21.800 41.800 22.200 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 0.600 13.100 1.000 13.500 ;
        RECT 11.800 12.800 12.200 13.200 ;
        RECT 16.600 18.800 17.000 19.200 ;
        RECT 15.800 14.800 16.200 15.200 ;
        RECT 10.200 11.800 10.600 12.200 ;
        RECT 15.800 12.800 16.200 13.200 ;
        RECT 22.200 16.800 22.600 17.200 ;
        RECT 20.600 15.800 21.000 16.200 ;
        RECT 23.800 13.800 24.200 14.200 ;
        RECT 29.400 18.800 29.800 19.200 ;
        RECT 31.000 13.100 31.400 13.500 ;
        RECT 39.800 11.800 40.200 12.200 ;
        RECT 2.200 6.800 2.600 7.200 ;
        RECT 17.400 8.800 17.800 9.200 ;
        RECT 11.800 7.800 12.200 8.200 ;
        RECT 10.200 6.800 10.600 7.200 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 13.400 5.800 13.800 6.200 ;
        RECT 19.000 6.800 19.400 7.200 ;
        RECT 19.000 5.800 19.400 6.200 ;
        RECT 21.400 6.600 21.800 7.000 ;
        RECT 23.000 6.800 23.400 7.200 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 23.800 5.800 24.200 6.200 ;
        RECT 25.400 5.800 25.800 6.200 ;
        RECT 36.600 4.800 37.000 5.200 ;
      LAYER metal2 ;
        RECT 0.600 25.100 1.000 27.900 ;
        RECT 2.200 23.100 2.600 28.900 ;
        RECT 3.800 26.100 4.200 26.200 ;
        RECT 4.600 26.100 5.000 26.200 ;
        RECT 3.800 25.800 5.000 26.100 ;
        RECT 7.000 23.100 7.400 28.900 ;
        RECT 19.800 28.800 20.200 29.200 ;
        RECT 19.800 28.200 20.100 28.800 ;
        RECT 13.400 27.800 13.800 28.200 ;
        RECT 17.400 28.100 17.800 28.200 ;
        RECT 16.600 27.800 17.800 28.100 ;
        RECT 19.800 27.800 20.200 28.200 ;
        RECT 20.600 27.800 21.000 28.200 ;
        RECT 24.600 28.100 25.000 28.200 ;
        RECT 23.800 27.800 25.000 28.100 ;
        RECT 13.400 27.000 13.700 27.800 ;
        RECT 13.400 26.600 13.800 27.000 ;
        RECT 10.200 26.100 10.600 26.200 ;
        RECT 11.000 26.100 11.400 26.200 ;
        RECT 10.200 25.800 11.400 26.100 ;
        RECT 9.400 21.800 9.800 22.200 ;
        RECT 0.600 13.100 1.000 15.900 ;
        RECT 2.200 12.100 2.600 17.900 ;
        RECT 5.400 14.800 5.800 15.200 ;
        RECT 5.400 9.200 5.700 14.800 ;
        RECT 7.000 12.100 7.400 17.900 ;
        RECT 9.400 14.200 9.700 21.800 ;
        RECT 16.600 19.200 16.900 27.800 ;
        RECT 17.400 26.100 17.700 27.800 ;
        RECT 19.000 27.100 19.400 27.200 ;
        RECT 19.000 26.800 20.100 27.100 ;
        RECT 18.200 26.100 18.600 26.200 ;
        RECT 17.400 25.800 18.600 26.100 ;
        RECT 16.600 18.800 17.000 19.200 ;
        RECT 19.000 16.800 19.400 17.200 ;
        RECT 19.000 15.200 19.300 16.800 ;
        RECT 15.800 14.800 16.200 15.200 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 9.400 13.800 9.800 14.200 ;
        RECT 11.800 13.800 12.200 14.200 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 11.800 13.200 12.100 13.800 ;
        RECT 11.800 12.800 12.200 13.200 ;
        RECT 10.200 11.800 10.600 12.200 ;
        RECT 5.400 8.800 5.800 9.200 ;
        RECT 7.000 7.800 7.400 8.200 ;
        RECT 1.400 7.100 1.800 7.200 ;
        RECT 2.200 7.100 2.600 7.200 ;
        RECT 1.400 6.800 2.600 7.100 ;
        RECT 7.000 6.200 7.300 7.800 ;
        RECT 10.200 7.200 10.500 11.800 ;
        RECT 11.800 7.800 12.200 8.200 ;
        RECT 10.200 6.800 10.600 7.200 ;
        RECT 11.800 6.200 12.100 7.800 ;
        RECT 13.400 6.200 13.700 13.800 ;
        RECT 15.800 13.200 16.100 14.800 ;
        RECT 19.800 14.200 20.100 26.800 ;
        RECT 20.600 22.200 20.900 27.800 ;
        RECT 23.000 26.800 23.400 27.200 ;
        RECT 21.400 26.100 21.800 26.200 ;
        RECT 22.200 26.100 22.600 26.200 ;
        RECT 21.400 25.800 22.600 26.100 ;
        RECT 20.600 21.800 21.000 22.200 ;
        RECT 23.000 17.200 23.300 26.800 ;
        RECT 23.800 26.200 24.100 27.800 ;
        RECT 23.800 25.800 24.200 26.200 ;
        RECT 29.400 26.100 29.800 26.200 ;
        RECT 30.200 26.100 30.600 26.200 ;
        RECT 29.400 25.800 30.600 26.100 ;
        RECT 31.800 25.800 32.200 26.200 ;
        RECT 23.800 19.200 24.100 25.800 ;
        RECT 31.800 25.200 32.100 25.800 ;
        RECT 31.800 24.800 32.200 25.200 ;
        RECT 32.600 25.100 33.000 27.900 ;
        RECT 34.200 23.100 34.600 28.900 ;
        RECT 35.800 25.800 36.200 26.200 ;
        RECT 35.800 25.200 36.100 25.800 ;
        RECT 35.800 24.800 36.200 25.200 ;
        RECT 39.000 23.100 39.400 28.900 ;
        RECT 41.400 21.800 41.800 22.200 ;
        RECT 23.800 18.800 24.200 19.200 ;
        RECT 28.600 19.100 29.000 19.200 ;
        RECT 29.400 19.100 29.800 19.200 ;
        RECT 28.600 18.800 29.800 19.100 ;
        RECT 22.200 17.100 22.600 17.200 ;
        RECT 23.000 17.100 23.400 17.200 ;
        RECT 22.200 16.800 23.400 17.100 ;
        RECT 20.600 15.800 21.000 16.200 ;
        RECT 25.400 15.800 25.800 16.200 ;
        RECT 19.000 14.100 19.400 14.200 ;
        RECT 19.800 14.100 20.200 14.200 ;
        RECT 19.000 13.800 20.200 14.100 ;
        RECT 15.800 13.100 16.200 13.200 ;
        RECT 16.600 13.100 17.000 13.200 ;
        RECT 15.800 12.800 17.000 13.100 ;
        RECT 17.400 11.800 17.800 12.200 ;
        RECT 17.400 11.200 17.700 11.800 ;
        RECT 17.400 10.800 17.800 11.200 ;
        RECT 14.200 9.800 14.600 10.200 ;
        RECT 14.200 7.200 14.500 9.800 ;
        RECT 20.600 9.200 20.900 15.800 ;
        RECT 21.400 14.800 21.800 15.200 ;
        RECT 21.400 12.200 21.700 14.800 ;
        RECT 25.400 14.200 25.700 15.800 ;
        RECT 27.000 14.800 27.400 15.200 ;
        RECT 23.800 13.800 24.200 14.200 ;
        RECT 25.400 13.800 25.800 14.200 ;
        RECT 26.200 13.800 26.600 14.200 ;
        RECT 22.200 13.100 22.600 13.200 ;
        RECT 23.000 13.100 23.400 13.200 ;
        RECT 22.200 12.800 23.400 13.100 ;
        RECT 21.400 11.800 21.800 12.200 ;
        RECT 15.000 8.800 15.400 9.200 ;
        RECT 17.400 9.100 17.800 9.200 ;
        RECT 18.200 9.100 18.600 9.200 ;
        RECT 17.400 8.800 18.600 9.100 ;
        RECT 20.600 8.800 21.000 9.200 ;
        RECT 15.000 8.200 15.300 8.800 ;
        RECT 15.000 7.800 15.400 8.200 ;
        RECT 15.800 7.800 16.200 8.200 ;
        RECT 16.600 7.800 17.000 8.200 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 15.800 6.200 16.100 7.800 ;
        RECT 16.600 7.200 16.900 7.800 ;
        RECT 16.600 6.800 17.000 7.200 ;
        RECT 19.000 7.100 19.400 7.200 ;
        RECT 19.000 6.800 20.100 7.100 ;
        RECT 19.800 6.200 20.100 6.800 ;
        RECT 21.400 7.000 21.700 11.800 ;
        RECT 23.800 10.200 24.100 13.800 ;
        RECT 24.600 11.800 25.000 12.200 ;
        RECT 23.800 9.800 24.200 10.200 ;
        RECT 22.200 8.100 22.600 8.200 ;
        RECT 23.000 8.100 23.400 8.200 ;
        RECT 22.200 7.800 23.400 8.100 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 23.800 7.100 24.100 9.800 ;
        RECT 24.600 8.200 24.900 11.800 ;
        RECT 26.200 9.200 26.500 13.800 ;
        RECT 27.000 12.200 27.300 14.800 ;
        RECT 31.000 13.100 31.400 15.900 ;
        RECT 27.000 11.800 27.400 12.200 ;
        RECT 32.600 12.100 33.000 17.900 ;
        RECT 33.400 14.700 33.800 15.100 ;
        RECT 25.400 8.800 25.800 9.200 ;
        RECT 26.200 8.800 26.600 9.200 ;
        RECT 24.600 7.800 25.000 8.200 ;
        RECT 21.400 6.600 21.800 7.000 ;
        RECT 23.000 6.800 24.100 7.100 ;
        RECT 25.400 6.200 25.700 8.800 ;
        RECT 26.200 8.200 26.500 8.800 ;
        RECT 26.200 7.800 26.600 8.200 ;
        RECT 27.000 7.200 27.300 11.800 ;
        RECT 33.400 9.200 33.700 14.700 ;
        RECT 36.600 11.800 37.000 12.200 ;
        RECT 37.400 12.100 37.800 17.900 ;
        RECT 38.200 16.800 38.600 17.200 ;
        RECT 38.200 15.200 38.500 16.800 ;
        RECT 41.400 15.200 41.700 21.800 ;
        RECT 38.200 14.800 38.600 15.200 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 33.400 8.100 33.800 8.200 ;
        RECT 34.200 8.100 34.600 8.200 ;
        RECT 33.400 7.800 34.600 8.100 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 4.600 6.100 5.000 6.200 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 4.600 5.800 5.800 6.100 ;
        RECT 7.000 5.800 7.400 6.200 ;
        RECT 11.800 5.800 12.200 6.200 ;
        RECT 13.400 5.800 13.800 6.200 ;
        RECT 15.800 5.800 16.200 6.200 ;
        RECT 18.200 6.100 18.600 6.200 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 18.200 5.800 19.400 6.100 ;
        RECT 19.800 5.800 20.200 6.200 ;
        RECT 23.000 6.100 23.400 6.200 ;
        RECT 23.800 6.100 24.200 6.200 ;
        RECT 23.000 5.800 24.200 6.100 ;
        RECT 25.400 5.800 25.800 6.200 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 31.800 6.100 32.200 6.200 ;
        RECT 31.000 5.800 32.200 6.100 ;
        RECT 34.200 6.100 34.600 6.200 ;
        RECT 35.000 6.100 35.400 6.200 ;
        RECT 34.200 5.800 35.400 6.100 ;
        RECT 36.600 5.200 36.900 11.800 ;
        RECT 38.200 7.200 38.500 14.800 ;
        RECT 39.000 12.100 39.400 12.200 ;
        RECT 39.800 12.100 40.200 12.200 ;
        RECT 39.000 11.800 40.200 12.100 ;
        RECT 38.200 6.800 38.600 7.200 ;
        RECT 38.200 6.100 38.600 6.200 ;
        RECT 39.000 6.100 39.400 6.200 ;
        RECT 38.200 5.800 39.400 6.100 ;
        RECT 36.600 4.800 37.000 5.200 ;
      LAYER via2 ;
        RECT 4.600 25.800 5.000 26.200 ;
        RECT 23.000 16.800 23.400 17.200 ;
        RECT 16.600 12.800 17.000 13.200 ;
        RECT 23.000 12.800 23.400 13.200 ;
        RECT 18.200 8.800 18.600 9.200 ;
        RECT 5.400 5.800 5.800 6.200 ;
        RECT 35.000 5.800 35.400 6.200 ;
      LAYER metal3 ;
        RECT 19.800 28.800 20.200 29.200 ;
        RECT 13.400 28.100 13.800 28.200 ;
        RECT 19.800 28.100 20.100 28.800 ;
        RECT 13.400 27.800 20.100 28.100 ;
        RECT 4.600 26.100 5.000 26.200 ;
        RECT 10.200 26.100 10.600 26.200 ;
        RECT 4.600 25.800 10.600 26.100 ;
        RECT 21.400 26.100 21.800 26.200 ;
        RECT 29.400 26.100 29.800 26.200 ;
        RECT 21.400 25.800 29.800 26.100 ;
        RECT 31.800 25.800 36.100 26.100 ;
        RECT 31.800 25.200 32.100 25.800 ;
        RECT 35.800 25.200 36.100 25.800 ;
        RECT 31.800 24.800 32.200 25.200 ;
        RECT 35.800 24.800 36.200 25.200 ;
        RECT 20.600 21.800 21.000 22.200 ;
        RECT 20.600 21.200 20.900 21.800 ;
        RECT 20.600 20.800 21.000 21.200 ;
        RECT 23.800 19.100 24.200 19.200 ;
        RECT 28.600 19.100 29.000 19.200 ;
        RECT 23.800 18.800 29.000 19.100 ;
        RECT 19.000 17.100 19.400 17.200 ;
        RECT 23.000 17.100 23.400 17.200 ;
        RECT 38.200 17.100 38.600 17.200 ;
        RECT 19.000 16.800 38.600 17.100 ;
        RECT 38.200 15.100 38.600 15.200 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 38.200 14.800 41.800 15.100 ;
        RECT 9.400 14.100 9.800 14.200 ;
        RECT 11.800 14.100 12.200 14.200 ;
        RECT 19.000 14.100 19.400 14.200 ;
        RECT 25.400 14.100 25.800 14.200 ;
        RECT 9.400 13.800 25.800 14.100 ;
        RECT 16.600 13.100 17.000 13.200 ;
        RECT 23.000 13.100 23.400 13.200 ;
        RECT 16.600 12.800 23.400 13.100 ;
        RECT 21.400 12.100 21.800 12.200 ;
        RECT 27.000 12.100 27.400 12.200 ;
        RECT 36.600 12.100 37.000 12.200 ;
        RECT 39.000 12.100 39.400 12.200 ;
        RECT 21.400 11.800 39.400 12.100 ;
        RECT 17.400 11.100 17.800 11.200 ;
        RECT 19.000 11.100 19.400 11.200 ;
        RECT 17.400 10.800 19.400 11.100 ;
        RECT 14.200 10.100 14.600 10.200 ;
        RECT 23.800 10.100 24.200 10.200 ;
        RECT 14.200 9.800 24.200 10.100 ;
        RECT 15.000 8.800 15.400 9.200 ;
        RECT 18.200 9.100 18.600 9.200 ;
        RECT 20.600 9.100 21.000 9.200 ;
        RECT 25.400 9.100 25.800 9.200 ;
        RECT 26.200 9.100 26.600 9.200 ;
        RECT 17.400 8.800 26.600 9.100 ;
        RECT 7.000 8.100 7.400 8.200 ;
        RECT 15.000 8.100 15.300 8.800 ;
        RECT 7.000 7.800 15.300 8.100 ;
        RECT 15.800 8.100 16.200 8.200 ;
        RECT 20.600 8.100 21.000 8.200 ;
        RECT 22.200 8.100 22.600 8.200 ;
        RECT 15.800 7.800 22.600 8.100 ;
        RECT 24.600 8.100 25.000 8.200 ;
        RECT 33.400 8.100 33.800 8.200 ;
        RECT 24.600 7.800 33.800 8.100 ;
        RECT 1.400 7.100 1.800 7.200 ;
        RECT 16.600 7.100 17.000 7.200 ;
        RECT 1.400 6.800 17.000 7.100 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 15.800 6.100 16.200 6.200 ;
        RECT 4.600 5.800 16.200 6.100 ;
        RECT 18.200 6.100 18.600 6.200 ;
        RECT 19.000 6.100 19.400 6.200 ;
        RECT 18.200 5.800 19.400 6.100 ;
        RECT 23.000 6.100 23.400 6.200 ;
        RECT 31.000 6.100 31.400 6.200 ;
        RECT 23.000 5.800 31.400 6.100 ;
        RECT 35.000 6.100 35.400 6.200 ;
        RECT 38.200 6.100 38.600 6.200 ;
        RECT 35.000 5.800 38.600 6.100 ;
      LAYER via3 ;
        RECT 19.000 10.800 19.400 11.200 ;
        RECT 20.600 7.800 21.000 8.200 ;
        RECT 19.000 5.800 19.400 6.200 ;
      LAYER metal4 ;
        RECT 20.600 20.800 21.000 21.200 ;
        RECT 19.000 10.800 19.400 11.200 ;
        RECT 19.000 6.200 19.300 10.800 ;
        RECT 20.600 8.200 20.900 20.800 ;
        RECT 20.600 7.800 21.000 8.200 ;
        RECT 19.000 5.800 19.400 6.200 ;
  END
END Watchdog
END LIBRARY

